USE WORK.config_pack.ALL;

PACKAGE project_pack IS

END;
