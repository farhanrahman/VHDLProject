LIBRARY IEEE;
USE IEEE.numeric_std.ALL;
USE IEEE.std_logic_1164.ALL;

PACKAGE cl_utility IS
	CONSTANT x_size 	: INTEGER := 6;
	CONSTANT p_size 	: INTEGER := 4;
	CONSTANT a_size 	: INTEGER := 8;
END PACKAGE cl_utility;